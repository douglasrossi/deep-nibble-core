-- Accumulator component