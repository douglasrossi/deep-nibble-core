library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity romx is
  port (
    i_ADDR : in std_logic_vector(4 downto 0);
    o_DATA : out std_logic_vector(14 downto 0)
  );
end romx;

architecture rtl of romx is

  type t_ROM is array(31 downto 0) of std_logic_vector(14 downto 0);

  constant c_MEM : t_ROM := (
    "000000000000000",
    "111111111111111",
    "111111111111110",
    "111111111111100",
    "111111111111000",
    "111111111110000",
    "111111111100000",
    "111111111000000",
    "111111110000000",
    "111111100000000",
    "111111000000000",
    "111110000000000",
    "111100000000000",
    "111000000000000",
    "110000000000000",
    "100000000000000",
    "000000000000000",
    "000000000000001",
    "000000000000010",
    "000000000000100",
    "000000000001000",
    "000000000010000",
    "000000000100000",
    "000000001000000",
    "000000010000000",
    "000000100000000",
    "000001000000000",
    "000010000000000",
    "000100000000000",
    "001000000000000",
    "010000000000000",
    "100000000000000");

begin

  o_DATA <= c_MEM(to_integer(unsigned(i_ADDR)));

end rtl;